library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 
entity sort_alg is

  port (
    rst : in std_logic;
    clk      : in std_logic;
 
    -- Inputs
    ain_tvalid   : in  std_logic;
    ain_tready	 : in  std_logic;
    ain_tdata 	 : in  std_logic_vector(15 downto 0);
    ain_tlast    : in  std_logic;
 
    -- Outputs
   	aout_tvalid  : out std_logic;
    aout_tready  : out std_logic;
    aout_tdata   : out std_logic_vector(15 downto 0);
    aout_tlast   : out std_logic
    );
end sort_alg;
 
architecture rtl of sort_alg is
  -- Memory
  type data_array is array (0 to 1023) of std_logic_vector(15 downto 0); -- max number of transactions is 1024
  signal data, sort_data : data_array := (others => (others => '0'));
   -- States for FSM
  type state_type is (idle, collect, assign, compare, check, increment, valid, ready, drive_one, drive_two);
  signal curr_state, next_state: state_type;
  -- Local signals
  signal i, j, d, x: integer := 0; -- Increment integers
  signal count: integer range 0 to 1023; -- field for number of transactions
  signal tmp_i, tmp_j: std_logic_vector(15 downto 0); -- Signals for temp values of data(i) and data(i+1)
   
  begin
  
  	process(clk, rst) is 
    begin
    if(rst = '1') then
    	curr_state <= idle;
    elsif(rising_edge(clk)) then
    	curr_state <= next_state;
	if(((ain_tvalid = '1') and (ain_tready = '1')) and ain_tlast = '0') then
		data(count) <= ain_tdata;
	end if;
	elsif(ain_tlast = '1') then
		next
    end if;
    end process;
    
    process(curr_state, ain_tdata, ain_tvalid, ain_tready) is
    begin
    case curr_state is
    	when idle =>
    	    aout_tdata <= (others => '0');
            aout_tvalid <= '0';
            aout_tready <= '0';
            aout_tlast <= '0';
            count <= 0;
            i <= 0;
            j <= 0;
            d <= 0;
            data <= (others => (others => '0'));
            if((ain_tvalid = '1') and (ain_tready = '1'))then
            	next_state <= collect;
            else
            	next_state <= idle;
	        end if;
        when collect =>
        	data(count) <= ain_tdata;
        	count <= count + 1;
            if(ain_tlast = '1') then
            	next_state <= assign;
            else
            	next_state <= collect;
            end if;
    	when assign =>
    	   tmp_i <= data(i);
    	   tmp_j <= data(i+1);
           next_state <= compare;
        when compare =>
            if(tmp_i > tmp_j) then
                data(i+1) <= tmp_i;
                data(i) <= tmp_j;
                next_state <= increment;
            else
                next_state <= increment;
            end if;
        when increment =>
            if(j /= count-2) then
                i <= i+1;
                next_state <= check;
            else
                next_state <= valid;
            end if;
            if(i = count-2) then
                j <= j+1;
            end if;
        when check =>
                if(i = count-1) then
                    i <= 0;
                    next_state <= assign;
                else
                    next_state <= assign;
                end if;
        when valid =>
        	aout_tvalid <= '1';
        	next_state <= ready;
        when ready =>
            aout_tready <= '1';
            next_state <= drive_one;
        when drive_one =>
            if(d /= count-1) then
                aout_tdata <= data(d);
                d <= d + 1;
                next_state <= drive_two;
            else
                aout_tlast <= '1';
                aout_tdata <= data(d);
                d <= 0;
            end if;
        when drive_two =>
            if(d /= count - 1) then
                aout_tdata <= data(d);
                next_state <= drive_one;
                d <= d + 1;
            else
                aout_tlast <= '1';
                aout_tdata <= data(d);
                d <= 0;
            end if;
    end case;
	end process;
end rtl;
